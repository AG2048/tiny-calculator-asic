/*
 * Copyright (c) 2025 Andy Gong
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module alu #(
    parameter DATA_WIDTH = 16
)(
    input  wire                   clk,        // clock
    input  wire                   rst_n,      // reset_n - low to reset
    // Add other ports as needed
);

endmodule